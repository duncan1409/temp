`timescale 1ns/100ps

module tb_ha(
    reg a, b,
    wire s, co
    );

    initial
    begin

    end
endmodule
